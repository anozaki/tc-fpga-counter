module BCDto7 (clk, rst, Input, Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] Input;
  output  wire [7:0] Output;

  TC_Constant # (.UUID(64'd2012982166399743991 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3F)) Constant8_0 (.out(wire_1));
  TC_Constant # (.UUID(64'd2550573772667337786 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_1 (.out(wire_16));
  TC_Constant # (.UUID(64'd4549024494436009822 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h5B)) Constant8_2 (.out(wire_30));
  TC_Constant # (.UUID(64'd998525519921564464 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h4F)) Constant8_3 (.out(wire_33));
  TC_Constant # (.UUID(64'd3920369487393325663 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h66)) Constant8_4 (.out(wire_25));
  TC_Constant # (.UUID(64'd2625829009698045294 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6D)) Constant8_5 (.out(wire_31));
  TC_Constant # (.UUID(64'd2346762579660488270 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7D)) Constant8_6 (.out(wire_17));
  TC_Constant # (.UUID(64'd1214826348397713202 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7)) Constant8_7 (.out(wire_23));
  TC_Constant # (.UUID(64'd3945780884569511531 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7F)) Constant8_8 (.out(wire_18));
  TC_Constant # (.UUID(64'd3169506249167528819 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6F)) Constant8_9 (.out(wire_36));
  TC_Switch # (.UUID(64'd2854467264430396311 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_10 (.en(wire_21), .in(wire_1), .out(wire_4_15));
  TC_Switch # (.UUID(64'd126247464589079487 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_11 (.en(wire_3), .in(wire_16), .out(wire_4_14));
  TC_Switch # (.UUID(64'd4194459744329446433 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_12 (.en(wire_5), .in(wire_30), .out(wire_4_13));
  TC_Switch # (.UUID(64'd3660124659456897319 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_13 (.en(wire_9), .in(wire_33), .out(wire_4_12));
  TC_Switch # (.UUID(64'd3479249487495867866 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_14 (.en(wire_22), .in(wire_25), .out(wire_4_11));
  TC_Switch # (.UUID(64'd164546049510304774 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_15 (.en(wire_0), .in(wire_31), .out(wire_4_10));
  TC_Switch # (.UUID(64'd2133161769490666473 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_16 (.en(wire_2), .in(wire_17), .out(wire_4_9));
  TC_Switch # (.UUID(64'd4498169374277615616 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_17 (.en(wire_20), .in(wire_23), .out(wire_4_8));
  TC_Switch # (.UUID(64'd2937706117705165057 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_18 (.en(wire_6), .in(wire_18), .out(wire_4_7));
  TC_Switch # (.UUID(64'd1787036094388788502 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_19 (.en(wire_34), .in(wire_36), .out(wire_4_4));
  TC_Constant # (.UUID(64'd1658099532637375037 ^ UUID), .BIT_WIDTH(64'd16), .value(16'h1)) Constant16_20 (.out(wire_32));
  TC_Shl # (.UUID(64'd1795661260779519106 ^ UUID), .BIT_WIDTH(64'd16)) Shl16_21 (.in(wire_32), .shift(wire_10), .out(wire_19));
  TC_Splitter16 # (.UUID(64'd1356072116386225699 ^ UUID)) Splitter16_22 (.in(wire_19), .out0(wire_8), .out1(wire_26));
  TC_Splitter8 # (.UUID(64'd941651416773416086 ^ UUID)) Splitter8_23 (.in(wire_8), .out0(wire_21), .out1(wire_3), .out2(wire_5), .out3(wire_9), .out4(wire_22), .out5(wire_0), .out6(wire_2), .out7(wire_20));
  TC_Constant # (.UUID(64'd2002483232534341337 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h77)) Constant8_24 (.out(wire_37));
  TC_Switch # (.UUID(64'd2857413362360145057 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_25 (.en(wire_7), .in(wire_37), .out(wire_4_2));
  TC_Constant # (.UUID(64'd1979438313497359298 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7C)) Constant8_26 (.out(wire_14));
  TC_Switch # (.UUID(64'd2008681196177291765 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_27 (.en(wire_24), .in(wire_14), .out(wire_4_0));
  TC_Constant # (.UUID(64'd4362291580534408181 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h39)) Constant8_28 (.out(wire_29));
  TC_Switch # (.UUID(64'd1693553741424283868 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_29 (.en(wire_13), .in(wire_29), .out(wire_4_1));
  TC_Constant # (.UUID(64'd3111790414817250394 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h5E)) Constant8_30 (.out(wire_27));
  TC_Switch # (.UUID(64'd1855426466790438356 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_31 (.en(wire_15), .in(wire_27), .out(wire_4_3));
  TC_Constant # (.UUID(64'd3217659841156582673 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h79)) Constant8_32 (.out(wire_11));
  TC_Switch # (.UUID(64'd168556671159170895 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_33 (.en(wire_28), .in(wire_11), .out(wire_4_5));
  TC_Constant # (.UUID(64'd2364403389279870864 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h71)) Constant8_34 (.out(wire_35));
  TC_Switch # (.UUID(64'd3591925781053722332 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_35 (.en(wire_12), .in(wire_35), .out(wire_4_6));
  TC_Splitter8 # (.UUID(64'd2573582878409240661 ^ UUID)) Splitter8_36 (.in(wire_26), .out0(wire_6), .out1(wire_34), .out2(wire_7), .out3(wire_24), .out4(wire_13), .out5(wire_15), .out6(wire_28), .out7(wire_12));

  wire [0:0] wire_0;
  wire [7:0] wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [7:0] wire_4;
  wire [7:0] wire_4_0;
  wire [7:0] wire_4_1;
  wire [7:0] wire_4_2;
  wire [7:0] wire_4_3;
  wire [7:0] wire_4_4;
  wire [7:0] wire_4_5;
  wire [7:0] wire_4_6;
  wire [7:0] wire_4_7;
  wire [7:0] wire_4_8;
  wire [7:0] wire_4_9;
  wire [7:0] wire_4_10;
  wire [7:0] wire_4_11;
  wire [7:0] wire_4_12;
  wire [7:0] wire_4_13;
  wire [7:0] wire_4_14;
  wire [7:0] wire_4_15;
  assign wire_4 = wire_4_0|wire_4_1|wire_4_2|wire_4_3|wire_4_4|wire_4_5|wire_4_6|wire_4_7|wire_4_8|wire_4_9|wire_4_10|wire_4_11|wire_4_12|wire_4_13|wire_4_14|wire_4_15;
  assign Output = wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [7:0] wire_8;
  wire [0:0] wire_9;
  wire [7:0] wire_10;
  assign wire_10 = Input;
  wire [7:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [7:0] wire_14;
  wire [0:0] wire_15;
  wire [7:0] wire_16;
  wire [7:0] wire_17;
  wire [7:0] wire_18;
  wire [15:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [7:0] wire_23;
  wire [0:0] wire_24;
  wire [7:0] wire_25;
  wire [7:0] wire_26;
  wire [7:0] wire_27;
  wire [0:0] wire_28;
  wire [7:0] wire_29;
  wire [7:0] wire_30;
  wire [7:0] wire_31;
  wire [15:0] wire_32;
  wire [7:0] wire_33;
  wire [0:0] wire_34;
  wire [7:0] wire_35;
  wire [7:0] wire_36;
  wire [7:0] wire_37;

endmodule
