module BCDto7 (clk, rst, Input, Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] Input;
  output  wire [7:0] Output;

  TC_Constant # (.UUID(64'd2012982166399743991 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3F)) Constant8_0 (.out(wire_12));
  TC_Constant # (.UUID(64'd2550573772667337786 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_1 (.out(wire_11));
  TC_Constant # (.UUID(64'd4549024494436009822 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h5B)) Constant8_2 (.out(wire_20));
  TC_Constant # (.UUID(64'd998525519921564464 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h4F)) Constant8_3 (.out(wire_25));
  TC_Constant # (.UUID(64'd3920369487393325663 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h66)) Constant8_4 (.out(wire_18));
  TC_Constant # (.UUID(64'd2625829009698045294 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6D)) Constant8_5 (.out(wire_10));
  TC_Constant # (.UUID(64'd2346762579660488270 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7D)) Constant8_6 (.out(wire_24));
  TC_Constant # (.UUID(64'd1214826348397713202 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7)) Constant8_7 (.out(wire_16));
  TC_Constant # (.UUID(64'd3945780884569511531 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7F)) Constant8_8 (.out(wire_7));
  TC_Constant # (.UUID(64'd3169506249167528819 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6F)) Constant8_9 (.out(wire_19));
  TC_Switch # (.UUID(64'd2854467264430396311 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_10 (.en(wire_0), .in(wire_12), .out(wire_2_8));
  TC_Switch # (.UUID(64'd126247464589079487 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_11 (.en(wire_13), .in(wire_11), .out(wire_2_6));
  TC_Switch # (.UUID(64'd4194459744329446433 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_12 (.en(wire_5), .in(wire_20), .out(wire_2_4));
  TC_Switch # (.UUID(64'd3660124659456897319 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_13 (.en(wire_4), .in(wire_25), .out(wire_2_2));
  TC_Switch # (.UUID(64'd3479249487495867866 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_14 (.en(wire_6), .in(wire_18), .out(wire_2_0));
  TC_Switch # (.UUID(64'd164546049510304774 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_15 (.en(wire_9), .in(wire_10), .out(wire_2_1));
  TC_Switch # (.UUID(64'd2133161769490666473 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_16 (.en(wire_22), .in(wire_24), .out(wire_2_3));
  TC_Switch # (.UUID(64'd4498169374277615616 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_17 (.en(wire_8), .in(wire_16), .out(wire_2_5));
  TC_Switch # (.UUID(64'd2937706117705165057 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_18 (.en(wire_1), .in(wire_7), .out(wire_2_7));
  TC_Switch # (.UUID(64'd1787036094388788502 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_19 (.en(wire_15), .in(wire_19), .out(wire_2_9));
  TC_Constant # (.UUID(64'd1658099532637375037 ^ UUID), .BIT_WIDTH(64'd16), .value(16'h1)) Constant16_20 (.out(wire_14));
  TC_Shl # (.UUID(64'd1795661260779519106 ^ UUID), .BIT_WIDTH(64'd16)) Shl16_21 (.in(wire_14), .shift(wire_23), .out(wire_3));
  TC_Splitter16 # (.UUID(64'd1356072116386225699 ^ UUID)) Splitter16_22 (.in(wire_3), .out0(wire_17), .out1(wire_21));
  TC_Splitter8 # (.UUID(64'd941651416773416086 ^ UUID)) Splitter8_23 (.in(wire_17), .out0(wire_0), .out1(wire_13), .out2(wire_5), .out3(wire_4), .out4(wire_6), .out5(wire_9), .out6(wire_22), .out7(wire_8));
  TC_Splitter8 # (.UUID(64'd2573582878409240661 ^ UUID)) Splitter8_24 (.in(wire_21), .out0(wire_1), .out1(wire_15), .out2(), .out3(), .out4(), .out5(), .out6(), .out7());

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [7:0] wire_2;
  wire [7:0] wire_2_0;
  wire [7:0] wire_2_1;
  wire [7:0] wire_2_2;
  wire [7:0] wire_2_3;
  wire [7:0] wire_2_4;
  wire [7:0] wire_2_5;
  wire [7:0] wire_2_6;
  wire [7:0] wire_2_7;
  wire [7:0] wire_2_8;
  wire [7:0] wire_2_9;
  assign wire_2 = wire_2_0|wire_2_1|wire_2_2|wire_2_3|wire_2_4|wire_2_5|wire_2_6|wire_2_7|wire_2_8|wire_2_9;
  assign Output = wire_2;
  wire [15:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [7:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [7:0] wire_10;
  wire [7:0] wire_11;
  wire [7:0] wire_12;
  wire [0:0] wire_13;
  wire [15:0] wire_14;
  wire [0:0] wire_15;
  wire [7:0] wire_16;
  wire [7:0] wire_17;
  wire [7:0] wire_18;
  wire [7:0] wire_19;
  wire [7:0] wire_20;
  wire [7:0] wire_21;
  wire [0:0] wire_22;
  wire [7:0] wire_23;
  assign wire_23 = Input;
  wire [7:0] wire_24;
  wire [7:0] wire_25;

endmodule
