module Count (clk, rst, hex, cycle, segtiming, debug, sel1, sel2, sel4, sel3, seg);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [0:0] hex;
  input  wire [31:0] cycle;
  input  wire [7:0] segtiming;
  output  wire [0:0] debug;
  output  wire [0:0] sel1;
  output  wire [0:0] sel2;
  output  wire [0:0] sel4;
  output  wire [0:0] sel3;
  output  wire [7:0] seg;

  TC_Counter # (.UUID(64'd2825092236961754806 ^ UUID), .BIT_WIDTH(64'd32), .count(32'd1)) Counter32_0 (.clk(clk), .rst(rst), .save(wire_3), .in(wire_9), .out(wire_36));
  TC_Equal # (.UUID(64'd2815436595443163428 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_1 (.in0(wire_36), .in1(wire_18), .out(wire_3));
  TC_Constant # (.UUID(64'd2195057612476342464 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h0)) Constant32_2 (.out(wire_9));
  TC_Constant # (.UUID(64'd546252498989508678 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_3 (.out(wire_46));
  TC_Not # (.UUID(64'd2422787759609528762 ^ UUID), .BIT_WIDTH(64'd1)) Not_4 (.in(wire_29), .out(wire_49));
  TC_BitMemory # (.UUID(64'd1705741650994387132 ^ UUID)) BitMemory_5 (.clk(clk), .rst(rst), .save(wire_3), .in(wire_49), .out(wire_29));
  TC_Counter # (.UUID(64'd483971983369626439 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd1)) Counter8_6 (.clk(clk), .rst(rst), .save(wire_0), .in(wire_19), .out(wire_34));
  TC_Splitter8 # (.UUID(64'd4101664230818326465 ^ UUID)) Splitter8_7 (.in(wire_20), .out0(wire_17), .out1(wire_22), .out2(wire_23), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd3597258672609514624 ^ UUID)) Decoder3_8 (.dis(1'd0), .sel0(wire_17), .sel1(wire_22), .sel2(wire_23), .out0(wire_24), .out1(), .out2(wire_32), .out3(), .out4(wire_13), .out5(), .out6(wire_11), .out7());
  TC_Equal # (.UUID(64'd117864268316446527 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_9 (.in0(wire_47), .in1(wire_34), .out(wire_0));
  TC_Add # (.UUID(64'd1980091076031166279 ^ UUID), .BIT_WIDTH(64'd8)) Add8_10 (.in0(wire_20), .in1(wire_44), .ci(1'd0), .out(wire_2), .co());
  TC_Constant # (.UUID(64'd2518862973311040322 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h0)) Constant8_11 (.out(wire_19));
  TC_Register # (.UUID(64'd2081291577489777194 ^ UUID), .BIT_WIDTH(64'd8)) Register8_12 (.clk(clk), .rst(rst), .load(wire_35), .save(wire_0), .in(wire_15), .out(wire_20));
  TC_Constant # (.UUID(64'd153928343309100327 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_13 (.out(wire_44));
  TC_Constant # (.UUID(64'd1286628564572084475 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_14 (.out(wire_35));
  TC_Mux # (.UUID(64'd2948685002671300977 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_15 (.sel(wire_37), .in0(wire_2), .in1(wire_42), .out(wire_15));
  TC_Constant # (.UUID(64'd3545286715238984315 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h0)) Constant8_16 (.out(wire_42));
  TC_Constant # (.UUID(64'd4122733212507919227 ^ UUID), .BIT_WIDTH(64'd16), .value(16'h1)) Constant16_17 (.out(wire_45));
  TC_Register # (.UUID(64'd1625823934977110048 ^ UUID), .BIT_WIDTH(64'd16)) Register16_18 (.clk(clk), .rst(rst), .load(wire_46), .save(wire_3), .in(wire_31), .out(wire_25));
  TC_Add # (.UUID(64'd122654855124550273 ^ UUID), .BIT_WIDTH(64'd16)) Add16_19 (.in0(wire_45), .in1(wire_25), .ci(1'd0), .out(wire_31), .co());
  TC_Mul # (.UUID(64'd3153334337711300085 ^ UUID), .BIT_WIDTH(64'd16)) DivMod16_20 (.in0(wire_25), .in1(wire_12), .out0(wire_30), .out1(wire_38));
  TC_Mul # (.UUID(64'd1019817654100684335 ^ UUID), .BIT_WIDTH(64'd16)) DivMod16_21 (.in0(wire_30), .in1(wire_12), .out0(wire_14), .out1(wire_40));
  TC_Mul # (.UUID(64'd1272800169210062040 ^ UUID), .BIT_WIDTH(64'd16)) DivMod16_22 (.in0(wire_14), .in1(wire_12), .out0(wire_43), .out1(wire_33));
  TC_Mul # (.UUID(64'd2764462783378612215 ^ UUID), .BIT_WIDTH(64'd16)) DivMod16_23 (.in0(wire_43), .in1(wire_12), .out0(), .out1(wire_7));
  TC_Constant # (.UUID(64'd2381158419837267810 ^ UUID), .BIT_WIDTH(64'd16), .value(16'hA)) Constant16_24 (.out(wire_12));
  TC_Switch # (.UUID(64'd256255929719074981 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_25 (.en(wire_24), .in(wire_6), .out(wire_5_3));
  TC_Switch # (.UUID(64'd2563149550945562995 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_26 (.en(wire_32), .in(wire_27), .out(wire_5_2));
  TC_Switch # (.UUID(64'd581565553225179143 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_27 (.en(wire_13), .in(wire_26), .out(wire_5_1));
  TC_Switch # (.UUID(64'd737480421798412485 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_28 (.en(wire_11), .in(wire_28), .out(wire_5_0));
  TC_IndexerBit # (.UUID(64'd2496807660048089843 ^ UUID), .INDEX(64'd3)) IndexerBit_29 (.in({{56{1'b0}}, wire_2 }), .out(wire_37));
  TC_Shr # (.UUID(64'd998018581472987639 ^ UUID), .BIT_WIDTH(64'd16)) Shr16_30 (.in(wire_25), .shift(wire_8), .out(wire_1));
  TC_Mux # (.UUID(64'd3083196977234481570 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_31 (.sel(wire_4), .in0(wire_38[7:0]), .in1(wire_25[7:0]), .out(wire_16));
  TC_Mux # (.UUID(64'd4288529005240128355 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_32 (.sel(wire_4), .in0(wire_40[7:0]), .in1(wire_1[7:0]), .out(wire_50));
  TC_Mux # (.UUID(64'd711062639695075971 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_33 (.sel(wire_4), .in0(wire_33[7:0]), .in1(wire_10[7:0]), .out(wire_41));
  TC_Mux # (.UUID(64'd605319909683182157 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_34 (.sel(wire_4), .in0(wire_7[7:0]), .in1(wire_48[7:0]), .out(wire_39));
  TC_Shr # (.UUID(64'd3691018399315671673 ^ UUID), .BIT_WIDTH(64'd16)) Shr16_35 (.in(wire_1), .shift(wire_8), .out(wire_10));
  TC_Shr # (.UUID(64'd4051741116473833853 ^ UUID), .BIT_WIDTH(64'd16)) Shr16_36 (.in(wire_10), .shift(wire_8), .out(wire_48));
  TC_Constant # (.UUID(64'd3169403740848913423 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h4)) Constant8_37 (.out(wire_8));
  BCDto7 # (.UUID(64'd1597852324588432281 ^ UUID)) BCDto7_38 (.clk(clk), .rst(rst), .Input(wire_16), .Output(wire_6));
  BCDto7 # (.UUID(64'd2214513227759376550 ^ UUID)) BCDto7_39 (.clk(clk), .rst(rst), .Input(wire_50), .Output(wire_27));
  BCDto7 # (.UUID(64'd3044709782342299070 ^ UUID)) BCDto7_40 (.clk(clk), .rst(rst), .Input(wire_41), .Output(wire_26));
  BCDto7 # (.UUID(64'd1468960662727354083 ^ UUID)) BCDto7_41 (.clk(clk), .rst(rst), .Input(wire_39), .Output(wire_28));
  debounce # (.UUID(64'd2856614444045816445 ^ UUID)) debounce_42 (.clk(clk), .rst(rst), .Input(wire_21), .Output(wire_4));

  wire [0:0] wire_0;
  wire [15:0] wire_1;
  wire [7:0] wire_2;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [7:0] wire_5;
  wire [7:0] wire_5_0;
  wire [7:0] wire_5_1;
  wire [7:0] wire_5_2;
  wire [7:0] wire_5_3;
  assign wire_5 = wire_5_0|wire_5_1|wire_5_2|wire_5_3;
  assign seg = wire_5;
  wire [7:0] wire_6;
  wire [15:0] wire_7;
  wire [7:0] wire_8;
  wire [31:0] wire_9;
  wire [15:0] wire_10;
  wire [0:0] wire_11;
  assign sel4 = wire_11;
  wire [15:0] wire_12;
  wire [0:0] wire_13;
  assign sel3 = wire_13;
  wire [15:0] wire_14;
  wire [7:0] wire_15;
  wire [7:0] wire_16;
  wire [0:0] wire_17;
  wire [31:0] wire_18;
  assign wire_18 = cycle;
  wire [7:0] wire_19;
  wire [7:0] wire_20;
  wire [0:0] wire_21;
  assign wire_21 = hex;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  assign sel1 = wire_24;
  wire [15:0] wire_25;
  wire [7:0] wire_26;
  wire [7:0] wire_27;
  wire [7:0] wire_28;
  wire [0:0] wire_29;
  assign debug = wire_29;
  wire [15:0] wire_30;
  wire [15:0] wire_31;
  wire [0:0] wire_32;
  assign sel2 = wire_32;
  wire [15:0] wire_33;
  wire [7:0] wire_34;
  wire [0:0] wire_35;
  wire [31:0] wire_36;
  wire [0:0] wire_37;
  wire [15:0] wire_38;
  wire [7:0] wire_39;
  wire [15:0] wire_40;
  wire [7:0] wire_41;
  wire [7:0] wire_42;
  wire [15:0] wire_43;
  wire [7:0] wire_44;
  wire [15:0] wire_45;
  wire [0:0] wire_46;
  wire [7:0] wire_47;
  assign wire_47 = segtiming;
  wire [15:0] wire_48;
  wire [0:0] wire_49;
  wire [7:0] wire_50;

endmodule
