module Count (clk, rst, hex, cycle, segtiming, debug, sel1, sel2, sel4, sel3, seg);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [0:0] hex;
  input  wire [31:0] cycle;
  input  wire [7:0] segtiming;
  output  wire [0:0] debug;
  output  wire [0:0] sel1;
  output  wire [0:0] sel2;
  output  wire [0:0] sel4;
  output  wire [0:0] sel3;
  output  wire [7:0] seg;

  TC_Counter # (.UUID(64'd2825092236961754806 ^ UUID), .BIT_WIDTH(64'd32), .count(32'd1)) Counter32_0 (.clk(clk), .rst(rst), .save(wire_3), .in(wire_34), .out(wire_49));
  TC_Equal # (.UUID(64'd2815436595443163428 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_1 (.in0(wire_49), .in1(wire_38), .out(wire_3));
  TC_Constant # (.UUID(64'd2195057612476342464 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h0)) Constant32_2 (.out(wire_34));
  TC_Constant # (.UUID(64'd546252498989508678 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_3 (.out(wire_46));
  TC_Not # (.UUID(64'd2422787759609528762 ^ UUID), .BIT_WIDTH(64'd1)) Not_4 (.in(wire_35), .out(wire_21));
  TC_BitMemory # (.UUID(64'd1705741650994387132 ^ UUID)) BitMemory_5 (.clk(clk), .rst(rst), .save(wire_3), .in(wire_21), .out(wire_35));
  TC_Counter # (.UUID(64'd483971983369626439 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd1)) Counter8_6 (.clk(clk), .rst(rst), .save(wire_25), .in(wire_31), .out(wire_39));
  TC_Splitter8 # (.UUID(64'd4101664230818326465 ^ UUID)) Splitter8_7 (.in(wire_15), .out0(wire_41), .out1(wire_24), .out2(wire_17), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd3597258672609514624 ^ UUID)) Decoder3_8 (.dis(1'd0), .sel0(wire_41), .sel1(wire_24), .sel2(wire_17), .out0(wire_37), .out1(wire_6), .out2(wire_23), .out3(wire_4), .out4(), .out5(), .out6(), .out7());
  TC_Equal # (.UUID(64'd117864268316446527 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_9 (.in0(wire_26), .in1(wire_39), .out(wire_25));
  TC_Add # (.UUID(64'd1980091076031166279 ^ UUID), .BIT_WIDTH(64'd8)) Add8_10 (.in0(wire_15), .in1(wire_29), .ci(1'd0), .out(wire_16), .co());
  TC_Constant # (.UUID(64'd2518862973311040322 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h0)) Constant8_11 (.out(wire_31));
  TC_Register # (.UUID(64'd2081291577489777194 ^ UUID), .BIT_WIDTH(64'd8)) Register8_12 (.clk(clk), .rst(rst), .load(wire_40), .save(wire_25), .in(wire_0), .out(wire_15));
  TC_Constant # (.UUID(64'd153928343309100327 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_13 (.out(wire_29));
  TC_Constant # (.UUID(64'd1286628564572084475 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_14 (.out(wire_40));
  TC_Mux # (.UUID(64'd2948685002671300977 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_15 (.sel(wire_19), .in0(wire_16), .in1(wire_43), .out(wire_0));
  TC_Constant # (.UUID(64'd3545286715238984315 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h0)) Constant8_16 (.out(wire_43));
  TC_Constant # (.UUID(64'd4122733212507919227 ^ UUID), .BIT_WIDTH(64'd16), .value(16'h1)) Constant16_17 (.out(wire_18));
  TC_Register # (.UUID(64'd1625823934977110048 ^ UUID), .BIT_WIDTH(64'd16)) Register16_18 (.clk(clk), .rst(rst), .load(wire_46), .save(wire_3), .in(wire_7), .out(wire_13));
  TC_Add # (.UUID(64'd122654855124550273 ^ UUID), .BIT_WIDTH(64'd16)) Add16_19 (.in0(wire_18), .in1(wire_13), .ci(1'd0), .out(wire_7), .co());
  TC_Mul # (.UUID(64'd3153334337711300085 ^ UUID), .BIT_WIDTH(64'd16)) DivMod16_20 (.in0(wire_13), .in1(wire_14), .out0(wire_33), .out1(wire_32));
  TC_Mul # (.UUID(64'd1019817654100684335 ^ UUID), .BIT_WIDTH(64'd16)) DivMod16_21 (.in0(wire_33), .in1(wire_14), .out0(wire_30), .out1(wire_48));
  TC_Mul # (.UUID(64'd1272800169210062040 ^ UUID), .BIT_WIDTH(64'd16)) DivMod16_22 (.in0(wire_30), .in1(wire_14), .out0(wire_10), .out1(wire_45));
  TC_Mul # (.UUID(64'd2764462783378612215 ^ UUID), .BIT_WIDTH(64'd16)) DivMod16_23 (.in0(wire_10), .in1(wire_14), .out0(), .out1(wire_36));
  TC_Constant # (.UUID(64'd2381158419837267810 ^ UUID), .BIT_WIDTH(64'd16), .value(16'hA)) Constant16_24 (.out(wire_14));
  TC_Switch # (.UUID(64'd256255929719074981 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_25 (.en(wire_37), .in(wire_9), .out(wire_12_3));
  TC_Switch # (.UUID(64'd2563149550945562995 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_26 (.en(wire_6), .in(wire_8), .out(wire_12_2));
  TC_Switch # (.UUID(64'd581565553225179143 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_27 (.en(wire_23), .in(wire_1), .out(wire_12_1));
  TC_Switch # (.UUID(64'd737480421798412485 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_28 (.en(wire_4), .in(wire_22), .out(wire_12_0));
  TC_IndexerBit # (.UUID(64'd2496807660048089843 ^ UUID), .INDEX(64'd2)) IndexerBit_29 (.in({{56{1'b0}}, wire_16 }), .out(wire_19));
  TC_Shr # (.UUID(64'd998018581472987639 ^ UUID), .BIT_WIDTH(64'd16)) Shr16_30 (.in(wire_13), .shift(wire_5), .out(wire_28));
  TC_Mux # (.UUID(64'd3083196977234481570 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_31 (.sel(wire_2), .in0(wire_32[7:0]), .in1(wire_13[7:0]), .out(wire_42));
  TC_Mux # (.UUID(64'd4288529005240128355 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_32 (.sel(wire_2), .in0(wire_48[7:0]), .in1(wire_28[7:0]), .out(wire_27));
  TC_Mux # (.UUID(64'd711062639695075971 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_33 (.sel(wire_2), .in0(wire_45[7:0]), .in1(wire_11[7:0]), .out(wire_20));
  TC_Mux # (.UUID(64'd605319909683182157 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_34 (.sel(wire_2), .in0(wire_36[7:0]), .in1(wire_44[7:0]), .out(wire_47));
  TC_Shr # (.UUID(64'd3691018399315671673 ^ UUID), .BIT_WIDTH(64'd16)) Shr16_35 (.in(wire_28), .shift(wire_5), .out(wire_11));
  TC_Shr # (.UUID(64'd4051741116473833853 ^ UUID), .BIT_WIDTH(64'd16)) Shr16_36 (.in(wire_11), .shift(wire_5), .out(wire_44));
  BCDto7 # (.UUID(64'd1597852324588432281 ^ UUID)) BCDto7_37 (.clk(clk), .rst(rst), .Input(wire_42), .Output(wire_9));
  BCDto7 # (.UUID(64'd2214513227759376550 ^ UUID)) BCDto7_38 (.clk(clk), .rst(rst), .Input(wire_27), .Output(wire_8));
  BCDto7 # (.UUID(64'd3044709782342299070 ^ UUID)) BCDto7_39 (.clk(clk), .rst(rst), .Input(wire_20), .Output(wire_1));
  BCDto7 # (.UUID(64'd1468960662727354083 ^ UUID)) BCDto7_40 (.clk(clk), .rst(rst), .Input(wire_47), .Output(wire_22));
  TC_Constant # (.UUID(64'd3169403740848913423 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h4)) Constant8_41 (.out(wire_5));

  wire [7:0] wire_0;
  wire [7:0] wire_1;
  wire [0:0] wire_2;
  assign wire_2 = hex;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  assign sel4 = wire_4;
  wire [7:0] wire_5;
  wire [0:0] wire_6;
  assign sel2 = wire_6;
  wire [15:0] wire_7;
  wire [7:0] wire_8;
  wire [7:0] wire_9;
  wire [15:0] wire_10;
  wire [15:0] wire_11;
  wire [7:0] wire_12;
  wire [7:0] wire_12_0;
  wire [7:0] wire_12_1;
  wire [7:0] wire_12_2;
  wire [7:0] wire_12_3;
  assign wire_12 = wire_12_0|wire_12_1|wire_12_2|wire_12_3;
  assign seg = wire_12;
  wire [15:0] wire_13;
  wire [15:0] wire_14;
  wire [7:0] wire_15;
  wire [7:0] wire_16;
  wire [0:0] wire_17;
  wire [15:0] wire_18;
  wire [0:0] wire_19;
  wire [7:0] wire_20;
  wire [0:0] wire_21;
  wire [7:0] wire_22;
  wire [0:0] wire_23;
  assign sel3 = wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [7:0] wire_26;
  assign wire_26 = segtiming;
  wire [7:0] wire_27;
  wire [15:0] wire_28;
  wire [7:0] wire_29;
  wire [15:0] wire_30;
  wire [7:0] wire_31;
  wire [15:0] wire_32;
  wire [15:0] wire_33;
  wire [31:0] wire_34;
  wire [0:0] wire_35;
  assign debug = wire_35;
  wire [15:0] wire_36;
  wire [0:0] wire_37;
  assign sel1 = wire_37;
  wire [31:0] wire_38;
  assign wire_38 = cycle;
  wire [7:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [7:0] wire_42;
  wire [7:0] wire_43;
  wire [15:0] wire_44;
  wire [15:0] wire_45;
  wire [0:0] wire_46;
  wire [7:0] wire_47;
  wire [15:0] wire_48;
  wire [31:0] wire_49;

endmodule
